module register_file(
  input clk,
  input write_enable,
  input [2:0]read_reg1,
  input [2:0]read_reg2,
  input [2:0]write_reg,
  input [7:0]write_data,
  output [7:0]read_data1,
  output [7:0]read_data2);
  reg[7:0] registers[7:0];
  assign read_data1= registers[read_reg1];
  assign read_data2= registers[read_reg2];
  always @(posedge clk) begin 
    if(write_enable)
      registers[write_reg]<=write_data;
  end 
endmodule
